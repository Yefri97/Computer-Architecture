library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity InstructionMemory is
    Port ( address : in  STD_LOGIC_VECTOR (31 downto 0);
           rst : in  STD_LOGIC;
           dataOut : out  STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type rom_type is array (127 downto 0) of std_logic_vector (31 downto 0);
signal ROM : rom_type := (	"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000000000000000000000000000000", "00000000000000000000000000000000", 
									"00000001000000000000000000000000", "00000001000000000000000000000000", 
									"01111111111111111111111111011000", "10111100000100000010000000000010", 
									"10111000000100000010000000000010", "10001100000100000010000000000001", 
									"10001010000100000010000000000011", "10001000000100000010000000000010", 
									"10111010000100000010000000000000", "00000001000000000000000000000000", 
									"10000001110000110110000000000010", "10010100000100000000000000010111", 
									"10101110000000101000000000001000", "00000001000000000000000000000000", 
									"01111111111111111111111111000100", "10110010000100000000000000001001", 
									"10110000000100000000000000000110", "00000001000000000000000000000000", 
									"01111111111111111111111111010110", "10110110000100000010000000000010", 
									"10110100000100000000000000011100", "10010100000100000000000000010111", 
									"10101110000000101000000000001000", "00000001000000000000000000000000", 
									"01111111111111111111111111001110", "10110010000100000000000000001001", 
									"10110000000100000000000000000101", "00000001000000000000000000000000", 
									"01111111111111111111111111100000", "10110110000100000010000000000001", 
									"10110100000100000000000000011100", "10010100000100000000000000010111", 
									"10101110000000101000000000001000", "00000001000000000000000000000000", 
									"01111111111111111111111111011000", "10110010000100000000000000001001", 
									"10110000000100000000000000000100", "00000001000000000000000000000000", 
									"01111111111111111111111111101010", "10110110000100000010000000000000", 
									"10110100000100000000000000011100", "10010100000100000010000000000000", 
									"10011010000100000000000000001111", "00000001000000000000000000000000", 
									"10000001110000111010000000000010", "00000001000000000000000000000000", 
									"00000110101111111111111111111000", "10000000101001000100000000011011", 
									"10100010000100000000000000010111", "10101110000001000110000000000001", 
									"10010010000100000000000000001000", "00000001000000000000000000000000", 
									"01111111111111111111111111101010", "10110010000100000000000000011010", 
									"10110000000100000000000000001001", "00000001000000000000000000000000", 
									"00000010100000000000000000001100", "10000000101001000100000000011011", 
									"10010010000100000010000000000001", "10100010000100000010000000000000", 
									"10011100000100000000000000001111", "00000001000000000000000000000000", 
									"10000001110000111110000000000010", "00000001000000000000000000000000", 
									"00000110101111111111111111111011", "10000000101001000000000000011001", 
									"10100000000100000000000000010111", "10101110000001000010000000000001", 
									"10010000000100000000000000010111", "10101110000000100000000000011000", 
									"00000001000000000000000000000000", "00000010100000000000000000001001", 
									"10000000101001000000000000011001", "10010000000100000010000000000000", 
									"10100000000100000010000000000000", "00000001000000000000000000000000", 
									"01000000000000000000000001000100", "00000001000000000000000000000000");

begin

process (rst, rom, address)
begin
	if (rst = '1') then
		-- Resetear
	else
		dataOut <= ROM(conv_integer(address(6 downto 0)));
	end if;
end process;

end Behavioral;